module top_module (
    output out);

//assign out = 1'b0;
    
    always @(*) begin
        out = 1'b0;
    end
    
endmodule
